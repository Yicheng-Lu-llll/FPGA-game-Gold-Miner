// nios_system.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module nios_system (
		input  wire        clk_clk,                  //               clk.clk
		input  wire [31:0] is_new_game_start_export, // is_new_game_start.export
		output wire [31:0] keycode_export,           //           keycode.export
		output wire [31:0] keycode0_export,          //          keycode0.export
		output wire [31:0] keycode1_export,          //          keycode1.export
		output wire [31:0] keycode2_export,          //          keycode2.export
		output wire [1:0]  otg_hpi_address_export,   //   otg_hpi_address.export
		output wire        otg_hpi_cs_export,        //        otg_hpi_cs.export
		input  wire [15:0] otg_hpi_data_in_port,     //      otg_hpi_data.in_port
		output wire [15:0] otg_hpi_data_out_port,    //                  .out_port
		output wire        otg_hpi_r_export,         //         otg_hpi_r.export
		output wire        otg_hpi_reset_export,     //     otg_hpi_reset.export
		output wire        otg_hpi_w_export,         //         otg_hpi_w.export
		output wire [31:0] position0_export,         //         position0.export
		output wire [31:0] position1_export,         //         position1.export
		output wire [31:0] position10_export,        //        position10.export
		output wire [31:0] position11_export,        //        position11.export
		output wire [31:0] position12_export,        //        position12.export
		output wire [31:0] position13_export,        //        position13.export
		output wire [31:0] position14_export,        //        position14.export
		output wire [31:0] position15_export,        //        position15.export
		output wire [31:0] position16_export,        //        position16.export
		output wire [31:0] position17_export,        //        position17.export
		output wire [31:0] position18_export,        //        position18.export
		output wire [31:0] position19_export,        //        position19.export
		output wire [31:0] position2_export,         //         position2.export
		output wire [31:0] position20_export,        //        position20.export
		output wire [31:0] position21_export,        //        position21.export
		output wire [31:0] position22_export,        //        position22.export
		output wire [31:0] position23_export,        //        position23.export
		output wire [31:0] position24_export,        //        position24.export
		output wire [31:0] position25_export,        //        position25.export
		output wire [31:0] position26_export,        //        position26.export
		output wire [31:0] position27_export,        //        position27.export
		output wire [31:0] position28_export,        //        position28.export
		output wire [31:0] position29_export,        //        position29.export
		output wire [31:0] position3_export,         //         position3.export
		output wire [31:0] position30_export,        //        position30.export
		output wire [31:0] position31_export,        //        position31.export
		output wire [31:0] position32_export,        //        position32.export
		output wire [31:0] position33_export,        //        position33.export
		output wire [31:0] position34_export,        //        position34.export
		output wire [31:0] position35_export,        //        position35.export
		output wire [31:0] position36_export,        //        position36.export
		output wire [31:0] position4_export,         //         position4.export
		output wire [31:0] position5_export,         //         position5.export
		output wire [31:0] position6_export,         //         position6.export
		output wire [31:0] position7_export,         //         position7.export
		output wire [31:0] position8_export,         //         position8.export
		output wire [31:0] position9_export,         //         position9.export
		input  wire        reset_reset_n,            //             reset.reset_n
		output wire        sdram_clk_clk,            //         sdram_clk.clk
		output wire [12:0] sdram_wire_addr,          //        sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,            //                  .ba
		output wire        sdram_wire_cas_n,         //                  .cas_n
		output wire        sdram_wire_cke,           //                  .cke
		output wire        sdram_wire_cs_n,          //                  .cs_n
		inout  wire [31:0] sdram_wire_dq,            //                  .dq
		output wire [3:0]  sdram_wire_dqm,           //                  .dqm
		output wire        sdram_wire_ras_n,         //                  .ras_n
		output wire        sdram_wire_we_n           //                  .we_n
	);

	wire         sdram_pll_c0_clk;                                            // sdram_pll:c0 -> [mm_interconnect_0:sdram_pll_c0_clk, rst_controller_002:clk, sdram:clk]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [28:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [28:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_readdata;              // sdram_pll:readdata -> mm_interconnect_0:sdram_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_sdram_pll_pll_slave_address;               // mm_interconnect_0:sdram_pll_pll_slave_address -> sdram_pll:address
	wire         mm_interconnect_0_sdram_pll_pll_slave_read;                  // mm_interconnect_0:sdram_pll_pll_slave_read -> sdram_pll:read
	wire         mm_interconnect_0_sdram_pll_pll_slave_write;                 // mm_interconnect_0:sdram_pll_pll_slave_write -> sdram_pll:write
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_writedata;             // mm_interconnect_0:sdram_pll_pll_slave_writedata -> sdram_pll:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [1:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                       // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                         // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                      // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                          // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                             // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                       // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                    // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                            // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                        // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_keycode_s1_chipselect;                     // mm_interconnect_0:keycode_s1_chipselect -> keycode:chipselect
	wire  [31:0] mm_interconnect_0_keycode_s1_readdata;                       // keycode:readdata -> mm_interconnect_0:keycode_s1_readdata
	wire   [1:0] mm_interconnect_0_keycode_s1_address;                        // mm_interconnect_0:keycode_s1_address -> keycode:address
	wire         mm_interconnect_0_keycode_s1_write;                          // mm_interconnect_0:keycode_s1_write -> keycode:write_n
	wire  [31:0] mm_interconnect_0_keycode_s1_writedata;                      // mm_interconnect_0:keycode_s1_writedata -> keycode:writedata
	wire         mm_interconnect_0_otg_hpi_address_s1_chipselect;             // mm_interconnect_0:otg_hpi_address_s1_chipselect -> otg_hpi_address:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_readdata;               // otg_hpi_address:readdata -> mm_interconnect_0:otg_hpi_address_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_address_s1_address;                // mm_interconnect_0:otg_hpi_address_s1_address -> otg_hpi_address:address
	wire         mm_interconnect_0_otg_hpi_address_s1_write;                  // mm_interconnect_0:otg_hpi_address_s1_write -> otg_hpi_address:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_writedata;              // mm_interconnect_0:otg_hpi_address_s1_writedata -> otg_hpi_address:writedata
	wire         mm_interconnect_0_otg_hpi_data_s1_chipselect;                // mm_interconnect_0:otg_hpi_data_s1_chipselect -> otg_hpi_data:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_readdata;                  // otg_hpi_data:readdata -> mm_interconnect_0:otg_hpi_data_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_data_s1_address;                   // mm_interconnect_0:otg_hpi_data_s1_address -> otg_hpi_data:address
	wire         mm_interconnect_0_otg_hpi_data_s1_write;                     // mm_interconnect_0:otg_hpi_data_s1_write -> otg_hpi_data:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_writedata;                 // mm_interconnect_0:otg_hpi_data_s1_writedata -> otg_hpi_data:writedata
	wire         mm_interconnect_0_otg_hpi_r_s1_chipselect;                   // mm_interconnect_0:otg_hpi_r_s1_chipselect -> otg_hpi_r:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_readdata;                     // otg_hpi_r:readdata -> mm_interconnect_0:otg_hpi_r_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_r_s1_address;                      // mm_interconnect_0:otg_hpi_r_s1_address -> otg_hpi_r:address
	wire         mm_interconnect_0_otg_hpi_r_s1_write;                        // mm_interconnect_0:otg_hpi_r_s1_write -> otg_hpi_r:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_writedata;                    // mm_interconnect_0:otg_hpi_r_s1_writedata -> otg_hpi_r:writedata
	wire         mm_interconnect_0_otg_hpi_w_s1_chipselect;                   // mm_interconnect_0:otg_hpi_w_s1_chipselect -> otg_hpi_w:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_readdata;                     // otg_hpi_w:readdata -> mm_interconnect_0:otg_hpi_w_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_w_s1_address;                      // mm_interconnect_0:otg_hpi_w_s1_address -> otg_hpi_w:address
	wire         mm_interconnect_0_otg_hpi_w_s1_write;                        // mm_interconnect_0:otg_hpi_w_s1_write -> otg_hpi_w:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_writedata;                    // mm_interconnect_0:otg_hpi_w_s1_writedata -> otg_hpi_w:writedata
	wire         mm_interconnect_0_otg_hpi_cs_s1_chipselect;                  // mm_interconnect_0:otg_hpi_cs_s1_chipselect -> otg_hpi_cs:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_readdata;                    // otg_hpi_cs:readdata -> mm_interconnect_0:otg_hpi_cs_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_cs_s1_address;                     // mm_interconnect_0:otg_hpi_cs_s1_address -> otg_hpi_cs:address
	wire         mm_interconnect_0_otg_hpi_cs_s1_write;                       // mm_interconnect_0:otg_hpi_cs_s1_write -> otg_hpi_cs:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_writedata;                   // mm_interconnect_0:otg_hpi_cs_s1_writedata -> otg_hpi_cs:writedata
	wire         mm_interconnect_0_otg_hpi_reset_s1_chipselect;               // mm_interconnect_0:otg_hpi_reset_s1_chipselect -> otg_hpi_reset:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_reset_s1_readdata;                 // otg_hpi_reset:readdata -> mm_interconnect_0:otg_hpi_reset_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_reset_s1_address;                  // mm_interconnect_0:otg_hpi_reset_s1_address -> otg_hpi_reset:address
	wire         mm_interconnect_0_otg_hpi_reset_s1_write;                    // mm_interconnect_0:otg_hpi_reset_s1_write -> otg_hpi_reset:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_reset_s1_writedata;                // mm_interconnect_0:otg_hpi_reset_s1_writedata -> otg_hpi_reset:writedata
	wire         mm_interconnect_0_keycode_0_s1_chipselect;                   // mm_interconnect_0:keycode_0_s1_chipselect -> keycode_0:chipselect
	wire  [31:0] mm_interconnect_0_keycode_0_s1_readdata;                     // keycode_0:readdata -> mm_interconnect_0:keycode_0_s1_readdata
	wire   [1:0] mm_interconnect_0_keycode_0_s1_address;                      // mm_interconnect_0:keycode_0_s1_address -> keycode_0:address
	wire         mm_interconnect_0_keycode_0_s1_write;                        // mm_interconnect_0:keycode_0_s1_write -> keycode_0:write_n
	wire  [31:0] mm_interconnect_0_keycode_0_s1_writedata;                    // mm_interconnect_0:keycode_0_s1_writedata -> keycode_0:writedata
	wire         mm_interconnect_0_keycode_1_s1_chipselect;                   // mm_interconnect_0:keycode_1_s1_chipselect -> keycode_1:chipselect
	wire  [31:0] mm_interconnect_0_keycode_1_s1_readdata;                     // keycode_1:readdata -> mm_interconnect_0:keycode_1_s1_readdata
	wire   [1:0] mm_interconnect_0_keycode_1_s1_address;                      // mm_interconnect_0:keycode_1_s1_address -> keycode_1:address
	wire         mm_interconnect_0_keycode_1_s1_write;                        // mm_interconnect_0:keycode_1_s1_write -> keycode_1:write_n
	wire  [31:0] mm_interconnect_0_keycode_1_s1_writedata;                    // mm_interconnect_0:keycode_1_s1_writedata -> keycode_1:writedata
	wire         mm_interconnect_0_keycode_2_s1_chipselect;                   // mm_interconnect_0:keycode_2_s1_chipselect -> keycode_2:chipselect
	wire  [31:0] mm_interconnect_0_keycode_2_s1_readdata;                     // keycode_2:readdata -> mm_interconnect_0:keycode_2_s1_readdata
	wire   [1:0] mm_interconnect_0_keycode_2_s1_address;                      // mm_interconnect_0:keycode_2_s1_address -> keycode_2:address
	wire         mm_interconnect_0_keycode_2_s1_write;                        // mm_interconnect_0:keycode_2_s1_write -> keycode_2:write_n
	wire  [31:0] mm_interconnect_0_keycode_2_s1_writedata;                    // mm_interconnect_0:keycode_2_s1_writedata -> keycode_2:writedata
	wire         mm_interconnect_0_position_0_s1_chipselect;                  // mm_interconnect_0:position_0_s1_chipselect -> position_0:chipselect
	wire  [31:0] mm_interconnect_0_position_0_s1_readdata;                    // position_0:readdata -> mm_interconnect_0:position_0_s1_readdata
	wire   [1:0] mm_interconnect_0_position_0_s1_address;                     // mm_interconnect_0:position_0_s1_address -> position_0:address
	wire         mm_interconnect_0_position_0_s1_write;                       // mm_interconnect_0:position_0_s1_write -> position_0:write_n
	wire  [31:0] mm_interconnect_0_position_0_s1_writedata;                   // mm_interconnect_0:position_0_s1_writedata -> position_0:writedata
	wire         mm_interconnect_0_position_1_s1_chipselect;                  // mm_interconnect_0:position_1_s1_chipselect -> position_1:chipselect
	wire  [31:0] mm_interconnect_0_position_1_s1_readdata;                    // position_1:readdata -> mm_interconnect_0:position_1_s1_readdata
	wire   [1:0] mm_interconnect_0_position_1_s1_address;                     // mm_interconnect_0:position_1_s1_address -> position_1:address
	wire         mm_interconnect_0_position_1_s1_write;                       // mm_interconnect_0:position_1_s1_write -> position_1:write_n
	wire  [31:0] mm_interconnect_0_position_1_s1_writedata;                   // mm_interconnect_0:position_1_s1_writedata -> position_1:writedata
	wire         mm_interconnect_0_position_2_s1_chipselect;                  // mm_interconnect_0:position_2_s1_chipselect -> position_2:chipselect
	wire  [31:0] mm_interconnect_0_position_2_s1_readdata;                    // position_2:readdata -> mm_interconnect_0:position_2_s1_readdata
	wire   [1:0] mm_interconnect_0_position_2_s1_address;                     // mm_interconnect_0:position_2_s1_address -> position_2:address
	wire         mm_interconnect_0_position_2_s1_write;                       // mm_interconnect_0:position_2_s1_write -> position_2:write_n
	wire  [31:0] mm_interconnect_0_position_2_s1_writedata;                   // mm_interconnect_0:position_2_s1_writedata -> position_2:writedata
	wire         mm_interconnect_0_position_3_s1_chipselect;                  // mm_interconnect_0:position_3_s1_chipselect -> position_3:chipselect
	wire  [31:0] mm_interconnect_0_position_3_s1_readdata;                    // position_3:readdata -> mm_interconnect_0:position_3_s1_readdata
	wire   [1:0] mm_interconnect_0_position_3_s1_address;                     // mm_interconnect_0:position_3_s1_address -> position_3:address
	wire         mm_interconnect_0_position_3_s1_write;                       // mm_interconnect_0:position_3_s1_write -> position_3:write_n
	wire  [31:0] mm_interconnect_0_position_3_s1_writedata;                   // mm_interconnect_0:position_3_s1_writedata -> position_3:writedata
	wire         mm_interconnect_0_position_4_s1_chipselect;                  // mm_interconnect_0:position_4_s1_chipselect -> position_4:chipselect
	wire  [31:0] mm_interconnect_0_position_4_s1_readdata;                    // position_4:readdata -> mm_interconnect_0:position_4_s1_readdata
	wire   [1:0] mm_interconnect_0_position_4_s1_address;                     // mm_interconnect_0:position_4_s1_address -> position_4:address
	wire         mm_interconnect_0_position_4_s1_write;                       // mm_interconnect_0:position_4_s1_write -> position_4:write_n
	wire  [31:0] mm_interconnect_0_position_4_s1_writedata;                   // mm_interconnect_0:position_4_s1_writedata -> position_4:writedata
	wire         mm_interconnect_0_position_5_s1_chipselect;                  // mm_interconnect_0:position_5_s1_chipselect -> position_5:chipselect
	wire  [31:0] mm_interconnect_0_position_5_s1_readdata;                    // position_5:readdata -> mm_interconnect_0:position_5_s1_readdata
	wire   [1:0] mm_interconnect_0_position_5_s1_address;                     // mm_interconnect_0:position_5_s1_address -> position_5:address
	wire         mm_interconnect_0_position_5_s1_write;                       // mm_interconnect_0:position_5_s1_write -> position_5:write_n
	wire  [31:0] mm_interconnect_0_position_5_s1_writedata;                   // mm_interconnect_0:position_5_s1_writedata -> position_5:writedata
	wire         mm_interconnect_0_position_6_s1_chipselect;                  // mm_interconnect_0:position_6_s1_chipselect -> position_6:chipselect
	wire  [31:0] mm_interconnect_0_position_6_s1_readdata;                    // position_6:readdata -> mm_interconnect_0:position_6_s1_readdata
	wire   [1:0] mm_interconnect_0_position_6_s1_address;                     // mm_interconnect_0:position_6_s1_address -> position_6:address
	wire         mm_interconnect_0_position_6_s1_write;                       // mm_interconnect_0:position_6_s1_write -> position_6:write_n
	wire  [31:0] mm_interconnect_0_position_6_s1_writedata;                   // mm_interconnect_0:position_6_s1_writedata -> position_6:writedata
	wire         mm_interconnect_0_position_7_s1_chipselect;                  // mm_interconnect_0:position_7_s1_chipselect -> position_7:chipselect
	wire  [31:0] mm_interconnect_0_position_7_s1_readdata;                    // position_7:readdata -> mm_interconnect_0:position_7_s1_readdata
	wire   [1:0] mm_interconnect_0_position_7_s1_address;                     // mm_interconnect_0:position_7_s1_address -> position_7:address
	wire         mm_interconnect_0_position_7_s1_write;                       // mm_interconnect_0:position_7_s1_write -> position_7:write_n
	wire  [31:0] mm_interconnect_0_position_7_s1_writedata;                   // mm_interconnect_0:position_7_s1_writedata -> position_7:writedata
	wire         mm_interconnect_0_position_8_s1_chipselect;                  // mm_interconnect_0:position_8_s1_chipselect -> position_8:chipselect
	wire  [31:0] mm_interconnect_0_position_8_s1_readdata;                    // position_8:readdata -> mm_interconnect_0:position_8_s1_readdata
	wire   [1:0] mm_interconnect_0_position_8_s1_address;                     // mm_interconnect_0:position_8_s1_address -> position_8:address
	wire         mm_interconnect_0_position_8_s1_write;                       // mm_interconnect_0:position_8_s1_write -> position_8:write_n
	wire  [31:0] mm_interconnect_0_position_8_s1_writedata;                   // mm_interconnect_0:position_8_s1_writedata -> position_8:writedata
	wire         mm_interconnect_0_position_9_s1_chipselect;                  // mm_interconnect_0:position_9_s1_chipselect -> position_9:chipselect
	wire  [31:0] mm_interconnect_0_position_9_s1_readdata;                    // position_9:readdata -> mm_interconnect_0:position_9_s1_readdata
	wire   [1:0] mm_interconnect_0_position_9_s1_address;                     // mm_interconnect_0:position_9_s1_address -> position_9:address
	wire         mm_interconnect_0_position_9_s1_write;                       // mm_interconnect_0:position_9_s1_write -> position_9:write_n
	wire  [31:0] mm_interconnect_0_position_9_s1_writedata;                   // mm_interconnect_0:position_9_s1_writedata -> position_9:writedata
	wire         mm_interconnect_0_position_10_s1_chipselect;                 // mm_interconnect_0:position_10_s1_chipselect -> position_10:chipselect
	wire  [31:0] mm_interconnect_0_position_10_s1_readdata;                   // position_10:readdata -> mm_interconnect_0:position_10_s1_readdata
	wire   [1:0] mm_interconnect_0_position_10_s1_address;                    // mm_interconnect_0:position_10_s1_address -> position_10:address
	wire         mm_interconnect_0_position_10_s1_write;                      // mm_interconnect_0:position_10_s1_write -> position_10:write_n
	wire  [31:0] mm_interconnect_0_position_10_s1_writedata;                  // mm_interconnect_0:position_10_s1_writedata -> position_10:writedata
	wire         mm_interconnect_0_position_11_s1_chipselect;                 // mm_interconnect_0:position_11_s1_chipselect -> position_11:chipselect
	wire  [31:0] mm_interconnect_0_position_11_s1_readdata;                   // position_11:readdata -> mm_interconnect_0:position_11_s1_readdata
	wire   [1:0] mm_interconnect_0_position_11_s1_address;                    // mm_interconnect_0:position_11_s1_address -> position_11:address
	wire         mm_interconnect_0_position_11_s1_write;                      // mm_interconnect_0:position_11_s1_write -> position_11:write_n
	wire  [31:0] mm_interconnect_0_position_11_s1_writedata;                  // mm_interconnect_0:position_11_s1_writedata -> position_11:writedata
	wire         mm_interconnect_0_position_12_s1_chipselect;                 // mm_interconnect_0:position_12_s1_chipselect -> position_12:chipselect
	wire  [31:0] mm_interconnect_0_position_12_s1_readdata;                   // position_12:readdata -> mm_interconnect_0:position_12_s1_readdata
	wire   [1:0] mm_interconnect_0_position_12_s1_address;                    // mm_interconnect_0:position_12_s1_address -> position_12:address
	wire         mm_interconnect_0_position_12_s1_write;                      // mm_interconnect_0:position_12_s1_write -> position_12:write_n
	wire  [31:0] mm_interconnect_0_position_12_s1_writedata;                  // mm_interconnect_0:position_12_s1_writedata -> position_12:writedata
	wire         mm_interconnect_0_position_13_s1_chipselect;                 // mm_interconnect_0:position_13_s1_chipselect -> position_13:chipselect
	wire  [31:0] mm_interconnect_0_position_13_s1_readdata;                   // position_13:readdata -> mm_interconnect_0:position_13_s1_readdata
	wire   [1:0] mm_interconnect_0_position_13_s1_address;                    // mm_interconnect_0:position_13_s1_address -> position_13:address
	wire         mm_interconnect_0_position_13_s1_write;                      // mm_interconnect_0:position_13_s1_write -> position_13:write_n
	wire  [31:0] mm_interconnect_0_position_13_s1_writedata;                  // mm_interconnect_0:position_13_s1_writedata -> position_13:writedata
	wire         mm_interconnect_0_position_14_s1_chipselect;                 // mm_interconnect_0:position_14_s1_chipselect -> position_14:chipselect
	wire  [31:0] mm_interconnect_0_position_14_s1_readdata;                   // position_14:readdata -> mm_interconnect_0:position_14_s1_readdata
	wire   [1:0] mm_interconnect_0_position_14_s1_address;                    // mm_interconnect_0:position_14_s1_address -> position_14:address
	wire         mm_interconnect_0_position_14_s1_write;                      // mm_interconnect_0:position_14_s1_write -> position_14:write_n
	wire  [31:0] mm_interconnect_0_position_14_s1_writedata;                  // mm_interconnect_0:position_14_s1_writedata -> position_14:writedata
	wire         mm_interconnect_0_position_15_s1_chipselect;                 // mm_interconnect_0:position_15_s1_chipselect -> position_15:chipselect
	wire  [31:0] mm_interconnect_0_position_15_s1_readdata;                   // position_15:readdata -> mm_interconnect_0:position_15_s1_readdata
	wire   [1:0] mm_interconnect_0_position_15_s1_address;                    // mm_interconnect_0:position_15_s1_address -> position_15:address
	wire         mm_interconnect_0_position_15_s1_write;                      // mm_interconnect_0:position_15_s1_write -> position_15:write_n
	wire  [31:0] mm_interconnect_0_position_15_s1_writedata;                  // mm_interconnect_0:position_15_s1_writedata -> position_15:writedata
	wire         mm_interconnect_0_position_16_s1_chipselect;                 // mm_interconnect_0:position_16_s1_chipselect -> position_16:chipselect
	wire  [31:0] mm_interconnect_0_position_16_s1_readdata;                   // position_16:readdata -> mm_interconnect_0:position_16_s1_readdata
	wire   [1:0] mm_interconnect_0_position_16_s1_address;                    // mm_interconnect_0:position_16_s1_address -> position_16:address
	wire         mm_interconnect_0_position_16_s1_write;                      // mm_interconnect_0:position_16_s1_write -> position_16:write_n
	wire  [31:0] mm_interconnect_0_position_16_s1_writedata;                  // mm_interconnect_0:position_16_s1_writedata -> position_16:writedata
	wire         mm_interconnect_0_position_17_s1_chipselect;                 // mm_interconnect_0:position_17_s1_chipselect -> position_17:chipselect
	wire  [31:0] mm_interconnect_0_position_17_s1_readdata;                   // position_17:readdata -> mm_interconnect_0:position_17_s1_readdata
	wire   [1:0] mm_interconnect_0_position_17_s1_address;                    // mm_interconnect_0:position_17_s1_address -> position_17:address
	wire         mm_interconnect_0_position_17_s1_write;                      // mm_interconnect_0:position_17_s1_write -> position_17:write_n
	wire  [31:0] mm_interconnect_0_position_17_s1_writedata;                  // mm_interconnect_0:position_17_s1_writedata -> position_17:writedata
	wire         mm_interconnect_0_position_18_s1_chipselect;                 // mm_interconnect_0:position_18_s1_chipselect -> position_18:chipselect
	wire  [31:0] mm_interconnect_0_position_18_s1_readdata;                   // position_18:readdata -> mm_interconnect_0:position_18_s1_readdata
	wire   [1:0] mm_interconnect_0_position_18_s1_address;                    // mm_interconnect_0:position_18_s1_address -> position_18:address
	wire         mm_interconnect_0_position_18_s1_write;                      // mm_interconnect_0:position_18_s1_write -> position_18:write_n
	wire  [31:0] mm_interconnect_0_position_18_s1_writedata;                  // mm_interconnect_0:position_18_s1_writedata -> position_18:writedata
	wire         mm_interconnect_0_position_19_s1_chipselect;                 // mm_interconnect_0:position_19_s1_chipselect -> position_19:chipselect
	wire  [31:0] mm_interconnect_0_position_19_s1_readdata;                   // position_19:readdata -> mm_interconnect_0:position_19_s1_readdata
	wire   [1:0] mm_interconnect_0_position_19_s1_address;                    // mm_interconnect_0:position_19_s1_address -> position_19:address
	wire         mm_interconnect_0_position_19_s1_write;                      // mm_interconnect_0:position_19_s1_write -> position_19:write_n
	wire  [31:0] mm_interconnect_0_position_19_s1_writedata;                  // mm_interconnect_0:position_19_s1_writedata -> position_19:writedata
	wire         mm_interconnect_0_position_20_s1_chipselect;                 // mm_interconnect_0:position_20_s1_chipselect -> position_20:chipselect
	wire  [31:0] mm_interconnect_0_position_20_s1_readdata;                   // position_20:readdata -> mm_interconnect_0:position_20_s1_readdata
	wire   [1:0] mm_interconnect_0_position_20_s1_address;                    // mm_interconnect_0:position_20_s1_address -> position_20:address
	wire         mm_interconnect_0_position_20_s1_write;                      // mm_interconnect_0:position_20_s1_write -> position_20:write_n
	wire  [31:0] mm_interconnect_0_position_20_s1_writedata;                  // mm_interconnect_0:position_20_s1_writedata -> position_20:writedata
	wire  [31:0] mm_interconnect_0_is_new_game_start_s1_readdata;             // is_new_game_start:readdata -> mm_interconnect_0:is_new_game_start_s1_readdata
	wire   [1:0] mm_interconnect_0_is_new_game_start_s1_address;              // mm_interconnect_0:is_new_game_start_s1_address -> is_new_game_start:address
	wire         mm_interconnect_0_position_21_s1_chipselect;                 // mm_interconnect_0:position_21_s1_chipselect -> position_21:chipselect
	wire  [31:0] mm_interconnect_0_position_21_s1_readdata;                   // position_21:readdata -> mm_interconnect_0:position_21_s1_readdata
	wire   [1:0] mm_interconnect_0_position_21_s1_address;                    // mm_interconnect_0:position_21_s1_address -> position_21:address
	wire         mm_interconnect_0_position_21_s1_write;                      // mm_interconnect_0:position_21_s1_write -> position_21:write_n
	wire  [31:0] mm_interconnect_0_position_21_s1_writedata;                  // mm_interconnect_0:position_21_s1_writedata -> position_21:writedata
	wire         mm_interconnect_0_position_22_s1_chipselect;                 // mm_interconnect_0:position_22_s1_chipselect -> position_22:chipselect
	wire  [31:0] mm_interconnect_0_position_22_s1_readdata;                   // position_22:readdata -> mm_interconnect_0:position_22_s1_readdata
	wire   [1:0] mm_interconnect_0_position_22_s1_address;                    // mm_interconnect_0:position_22_s1_address -> position_22:address
	wire         mm_interconnect_0_position_22_s1_write;                      // mm_interconnect_0:position_22_s1_write -> position_22:write_n
	wire  [31:0] mm_interconnect_0_position_22_s1_writedata;                  // mm_interconnect_0:position_22_s1_writedata -> position_22:writedata
	wire         mm_interconnect_0_position_23_s1_chipselect;                 // mm_interconnect_0:position_23_s1_chipselect -> position_23:chipselect
	wire  [31:0] mm_interconnect_0_position_23_s1_readdata;                   // position_23:readdata -> mm_interconnect_0:position_23_s1_readdata
	wire   [1:0] mm_interconnect_0_position_23_s1_address;                    // mm_interconnect_0:position_23_s1_address -> position_23:address
	wire         mm_interconnect_0_position_23_s1_write;                      // mm_interconnect_0:position_23_s1_write -> position_23:write_n
	wire  [31:0] mm_interconnect_0_position_23_s1_writedata;                  // mm_interconnect_0:position_23_s1_writedata -> position_23:writedata
	wire         mm_interconnect_0_position_24_s1_chipselect;                 // mm_interconnect_0:position_24_s1_chipselect -> position_24:chipselect
	wire  [31:0] mm_interconnect_0_position_24_s1_readdata;                   // position_24:readdata -> mm_interconnect_0:position_24_s1_readdata
	wire   [1:0] mm_interconnect_0_position_24_s1_address;                    // mm_interconnect_0:position_24_s1_address -> position_24:address
	wire         mm_interconnect_0_position_24_s1_write;                      // mm_interconnect_0:position_24_s1_write -> position_24:write_n
	wire  [31:0] mm_interconnect_0_position_24_s1_writedata;                  // mm_interconnect_0:position_24_s1_writedata -> position_24:writedata
	wire         mm_interconnect_0_position_25_s1_chipselect;                 // mm_interconnect_0:position_25_s1_chipselect -> position_25:chipselect
	wire  [31:0] mm_interconnect_0_position_25_s1_readdata;                   // position_25:readdata -> mm_interconnect_0:position_25_s1_readdata
	wire   [1:0] mm_interconnect_0_position_25_s1_address;                    // mm_interconnect_0:position_25_s1_address -> position_25:address
	wire         mm_interconnect_0_position_25_s1_write;                      // mm_interconnect_0:position_25_s1_write -> position_25:write_n
	wire  [31:0] mm_interconnect_0_position_25_s1_writedata;                  // mm_interconnect_0:position_25_s1_writedata -> position_25:writedata
	wire         mm_interconnect_0_position_26_s1_chipselect;                 // mm_interconnect_0:position_26_s1_chipselect -> position_26:chipselect
	wire  [31:0] mm_interconnect_0_position_26_s1_readdata;                   // position_26:readdata -> mm_interconnect_0:position_26_s1_readdata
	wire   [1:0] mm_interconnect_0_position_26_s1_address;                    // mm_interconnect_0:position_26_s1_address -> position_26:address
	wire         mm_interconnect_0_position_26_s1_write;                      // mm_interconnect_0:position_26_s1_write -> position_26:write_n
	wire  [31:0] mm_interconnect_0_position_26_s1_writedata;                  // mm_interconnect_0:position_26_s1_writedata -> position_26:writedata
	wire         mm_interconnect_0_position_27_s1_chipselect;                 // mm_interconnect_0:position_27_s1_chipselect -> position_27:chipselect
	wire  [31:0] mm_interconnect_0_position_27_s1_readdata;                   // position_27:readdata -> mm_interconnect_0:position_27_s1_readdata
	wire   [1:0] mm_interconnect_0_position_27_s1_address;                    // mm_interconnect_0:position_27_s1_address -> position_27:address
	wire         mm_interconnect_0_position_27_s1_write;                      // mm_interconnect_0:position_27_s1_write -> position_27:write_n
	wire  [31:0] mm_interconnect_0_position_27_s1_writedata;                  // mm_interconnect_0:position_27_s1_writedata -> position_27:writedata
	wire         mm_interconnect_0_position_28_s1_chipselect;                 // mm_interconnect_0:position_28_s1_chipselect -> position_28:chipselect
	wire  [31:0] mm_interconnect_0_position_28_s1_readdata;                   // position_28:readdata -> mm_interconnect_0:position_28_s1_readdata
	wire   [1:0] mm_interconnect_0_position_28_s1_address;                    // mm_interconnect_0:position_28_s1_address -> position_28:address
	wire         mm_interconnect_0_position_28_s1_write;                      // mm_interconnect_0:position_28_s1_write -> position_28:write_n
	wire  [31:0] mm_interconnect_0_position_28_s1_writedata;                  // mm_interconnect_0:position_28_s1_writedata -> position_28:writedata
	wire         mm_interconnect_0_position_29_s1_chipselect;                 // mm_interconnect_0:position_29_s1_chipselect -> position_29:chipselect
	wire  [31:0] mm_interconnect_0_position_29_s1_readdata;                   // position_29:readdata -> mm_interconnect_0:position_29_s1_readdata
	wire   [1:0] mm_interconnect_0_position_29_s1_address;                    // mm_interconnect_0:position_29_s1_address -> position_29:address
	wire         mm_interconnect_0_position_29_s1_write;                      // mm_interconnect_0:position_29_s1_write -> position_29:write_n
	wire  [31:0] mm_interconnect_0_position_29_s1_writedata;                  // mm_interconnect_0:position_29_s1_writedata -> position_29:writedata
	wire         mm_interconnect_0_position_30_s1_chipselect;                 // mm_interconnect_0:position_30_s1_chipselect -> position_30:chipselect
	wire  [31:0] mm_interconnect_0_position_30_s1_readdata;                   // position_30:readdata -> mm_interconnect_0:position_30_s1_readdata
	wire   [1:0] mm_interconnect_0_position_30_s1_address;                    // mm_interconnect_0:position_30_s1_address -> position_30:address
	wire         mm_interconnect_0_position_30_s1_write;                      // mm_interconnect_0:position_30_s1_write -> position_30:write_n
	wire  [31:0] mm_interconnect_0_position_30_s1_writedata;                  // mm_interconnect_0:position_30_s1_writedata -> position_30:writedata
	wire         mm_interconnect_0_position_31_s1_chipselect;                 // mm_interconnect_0:position_31_s1_chipselect -> position_31:chipselect
	wire  [31:0] mm_interconnect_0_position_31_s1_readdata;                   // position_31:readdata -> mm_interconnect_0:position_31_s1_readdata
	wire   [1:0] mm_interconnect_0_position_31_s1_address;                    // mm_interconnect_0:position_31_s1_address -> position_31:address
	wire         mm_interconnect_0_position_31_s1_write;                      // mm_interconnect_0:position_31_s1_write -> position_31:write_n
	wire  [31:0] mm_interconnect_0_position_31_s1_writedata;                  // mm_interconnect_0:position_31_s1_writedata -> position_31:writedata
	wire         mm_interconnect_0_position_32_s1_chipselect;                 // mm_interconnect_0:position_32_s1_chipselect -> position_32:chipselect
	wire  [31:0] mm_interconnect_0_position_32_s1_readdata;                   // position_32:readdata -> mm_interconnect_0:position_32_s1_readdata
	wire   [1:0] mm_interconnect_0_position_32_s1_address;                    // mm_interconnect_0:position_32_s1_address -> position_32:address
	wire         mm_interconnect_0_position_32_s1_write;                      // mm_interconnect_0:position_32_s1_write -> position_32:write_n
	wire  [31:0] mm_interconnect_0_position_32_s1_writedata;                  // mm_interconnect_0:position_32_s1_writedata -> position_32:writedata
	wire         mm_interconnect_0_position_33_s1_chipselect;                 // mm_interconnect_0:position_33_s1_chipselect -> position_33:chipselect
	wire  [31:0] mm_interconnect_0_position_33_s1_readdata;                   // position_33:readdata -> mm_interconnect_0:position_33_s1_readdata
	wire   [1:0] mm_interconnect_0_position_33_s1_address;                    // mm_interconnect_0:position_33_s1_address -> position_33:address
	wire         mm_interconnect_0_position_33_s1_write;                      // mm_interconnect_0:position_33_s1_write -> position_33:write_n
	wire  [31:0] mm_interconnect_0_position_33_s1_writedata;                  // mm_interconnect_0:position_33_s1_writedata -> position_33:writedata
	wire         mm_interconnect_0_position_34_s1_chipselect;                 // mm_interconnect_0:position_34_s1_chipselect -> position_34:chipselect
	wire  [31:0] mm_interconnect_0_position_34_s1_readdata;                   // position_34:readdata -> mm_interconnect_0:position_34_s1_readdata
	wire   [1:0] mm_interconnect_0_position_34_s1_address;                    // mm_interconnect_0:position_34_s1_address -> position_34:address
	wire         mm_interconnect_0_position_34_s1_write;                      // mm_interconnect_0:position_34_s1_write -> position_34:write_n
	wire  [31:0] mm_interconnect_0_position_34_s1_writedata;                  // mm_interconnect_0:position_34_s1_writedata -> position_34:writedata
	wire         mm_interconnect_0_position_35_s1_chipselect;                 // mm_interconnect_0:position_35_s1_chipselect -> position_35:chipselect
	wire  [31:0] mm_interconnect_0_position_35_s1_readdata;                   // position_35:readdata -> mm_interconnect_0:position_35_s1_readdata
	wire   [1:0] mm_interconnect_0_position_35_s1_address;                    // mm_interconnect_0:position_35_s1_address -> position_35:address
	wire         mm_interconnect_0_position_35_s1_write;                      // mm_interconnect_0:position_35_s1_write -> position_35:write_n
	wire  [31:0] mm_interconnect_0_position_35_s1_writedata;                  // mm_interconnect_0:position_35_s1_writedata -> position_35:writedata
	wire         mm_interconnect_0_position_36_s1_chipselect;                 // mm_interconnect_0:position_36_s1_chipselect -> position_36:chipselect
	wire  [31:0] mm_interconnect_0_position_36_s1_readdata;                   // position_36:readdata -> mm_interconnect_0:position_36_s1_readdata
	wire   [1:0] mm_interconnect_0_position_36_s1_address;                    // mm_interconnect_0:position_36_s1_address -> position_36:address
	wire         mm_interconnect_0_position_36_s1_write;                      // mm_interconnect_0:position_36_s1_write -> position_36:write_n
	wire  [31:0] mm_interconnect_0_position_36_s1_writedata;                  // mm_interconnect_0:position_36_s1_writedata -> position_36:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [is_new_game_start:reset_n, jtag_uart_0:rst_n, keycode:reset_n, keycode_0:reset_n, keycode_1:reset_n, keycode_2:reset_n, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, otg_hpi_address:reset_n, otg_hpi_cs:reset_n, otg_hpi_data:reset_n, otg_hpi_r:reset_n, otg_hpi_reset:reset_n, otg_hpi_w:reset_n, position_0:reset_n, position_10:reset_n, position_11:reset_n, position_12:reset_n, position_13:reset_n, position_14:reset_n, position_15:reset_n, position_16:reset_n, position_17:reset_n, position_18:reset_n, position_19:reset_n, position_1:reset_n, position_20:reset_n, position_21:reset_n, position_22:reset_n, position_23:reset_n, position_24:reset_n, position_25:reset_n, position_26:reset_n, position_27:reset_n, position_28:reset_n, position_29:reset_n, position_2:reset_n, position_30:reset_n, position_31:reset_n, position_32:reset_n, position_33:reset_n, position_34:reset_n, position_35:reset_n, position_36:reset_n, position_3:reset_n, position_4:reset_n, position_5:reset_n, position_6:reset_n, position_7:reset_n, position_8:reset_n, position_9:reset_n]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, sdram_pll:reset, sysid_qsys_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_002_reset_out_reset;                          // rst_controller_002:reset_out -> [mm_interconnect_0:sdram_reset_reset_bridge_in_reset_reset, sdram:reset_n]

	nios_system_is_new_game_start is_new_game_start (
		.clk      (clk_clk),                                         //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address  (mm_interconnect_0_is_new_game_start_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_is_new_game_start_s1_readdata), //                    .readdata
		.in_port  (is_new_game_start_export)                         // external_connection.export
	);

	nios_system_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios_system_keycode keycode (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_keycode_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keycode_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keycode_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keycode_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keycode_s1_readdata),   //                    .readdata
		.out_port   (keycode_export)                           // external_connection.export
	);

	nios_system_keycode keycode_0 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_keycode_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keycode_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keycode_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keycode_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keycode_0_s1_readdata),   //                    .readdata
		.out_port   (keycode0_export)                            // external_connection.export
	);

	nios_system_keycode keycode_1 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_keycode_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keycode_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keycode_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keycode_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keycode_1_s1_readdata),   //                    .readdata
		.out_port   (keycode1_export)                            // external_connection.export
	);

	nios_system_keycode keycode_2 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_keycode_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keycode_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keycode_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keycode_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keycode_2_s1_readdata),   //                    .readdata
		.out_port   (keycode2_export)                            // external_connection.export
	);

	nios_system_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	nios_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	nios_system_otg_hpi_address otg_hpi_address (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_address_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_address_export)                           // external_connection.export
	);

	nios_system_otg_hpi_cs otg_hpi_cs (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_cs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_cs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_cs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_cs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_cs_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_cs_export)                           // external_connection.export
	);

	nios_system_otg_hpi_data otg_hpi_data (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_data_s1_readdata),   //                    .readdata
		.in_port    (otg_hpi_data_in_port),                         // external_connection.export
		.out_port   (otg_hpi_data_out_port)                         //                    .export
	);

	nios_system_otg_hpi_cs otg_hpi_r (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_r_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_r_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_r_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_r_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_r_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_r_export)                           // external_connection.export
	);

	nios_system_otg_hpi_cs otg_hpi_reset (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_reset_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_reset_export)                           // external_connection.export
	);

	nios_system_otg_hpi_cs otg_hpi_w (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_w_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_w_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_w_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_w_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_w_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_w_export)                           // external_connection.export
	);

	nios_system_keycode position_0 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_position_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_0_s1_readdata),   //                    .readdata
		.out_port   (position0_export)                            // external_connection.export
	);

	nios_system_keycode position_1 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_position_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_1_s1_readdata),   //                    .readdata
		.out_port   (position1_export)                            // external_connection.export
	);

	nios_system_keycode position_10 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_10_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_10_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_10_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_10_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_10_s1_readdata),   //                    .readdata
		.out_port   (position10_export)                            // external_connection.export
	);

	nios_system_keycode position_11 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_11_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_11_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_11_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_11_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_11_s1_readdata),   //                    .readdata
		.out_port   (position11_export)                            // external_connection.export
	);

	nios_system_keycode position_12 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_12_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_12_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_12_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_12_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_12_s1_readdata),   //                    .readdata
		.out_port   (position12_export)                            // external_connection.export
	);

	nios_system_keycode position_13 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_13_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_13_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_13_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_13_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_13_s1_readdata),   //                    .readdata
		.out_port   (position13_export)                            // external_connection.export
	);

	nios_system_keycode position_14 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_14_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_14_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_14_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_14_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_14_s1_readdata),   //                    .readdata
		.out_port   (position14_export)                            // external_connection.export
	);

	nios_system_keycode position_15 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_15_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_15_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_15_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_15_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_15_s1_readdata),   //                    .readdata
		.out_port   (position15_export)                            // external_connection.export
	);

	nios_system_keycode position_16 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_16_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_16_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_16_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_16_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_16_s1_readdata),   //                    .readdata
		.out_port   (position16_export)                            // external_connection.export
	);

	nios_system_keycode position_17 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_17_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_17_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_17_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_17_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_17_s1_readdata),   //                    .readdata
		.out_port   (position17_export)                            // external_connection.export
	);

	nios_system_keycode position_18 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_18_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_18_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_18_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_18_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_18_s1_readdata),   //                    .readdata
		.out_port   (position18_export)                            // external_connection.export
	);

	nios_system_keycode position_19 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_19_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_19_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_19_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_19_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_19_s1_readdata),   //                    .readdata
		.out_port   (position19_export)                            // external_connection.export
	);

	nios_system_keycode position_2 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_position_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_2_s1_readdata),   //                    .readdata
		.out_port   (position2_export)                            // external_connection.export
	);

	nios_system_keycode position_20 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_20_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_20_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_20_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_20_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_20_s1_readdata),   //                    .readdata
		.out_port   (position20_export)                            // external_connection.export
	);

	nios_system_keycode position_21 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_21_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_21_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_21_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_21_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_21_s1_readdata),   //                    .readdata
		.out_port   (position21_export)                            // external_connection.export
	);

	nios_system_keycode position_22 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_22_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_22_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_22_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_22_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_22_s1_readdata),   //                    .readdata
		.out_port   (position22_export)                            // external_connection.export
	);

	nios_system_keycode position_23 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_23_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_23_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_23_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_23_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_23_s1_readdata),   //                    .readdata
		.out_port   (position23_export)                            // external_connection.export
	);

	nios_system_keycode position_24 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_24_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_24_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_24_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_24_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_24_s1_readdata),   //                    .readdata
		.out_port   (position24_export)                            // external_connection.export
	);

	nios_system_keycode position_25 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_25_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_25_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_25_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_25_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_25_s1_readdata),   //                    .readdata
		.out_port   (position25_export)                            // external_connection.export
	);

	nios_system_keycode position_26 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_26_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_26_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_26_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_26_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_26_s1_readdata),   //                    .readdata
		.out_port   (position26_export)                            // external_connection.export
	);

	nios_system_keycode position_27 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_27_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_27_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_27_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_27_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_27_s1_readdata),   //                    .readdata
		.out_port   (position27_export)                            // external_connection.export
	);

	nios_system_keycode position_28 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_28_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_28_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_28_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_28_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_28_s1_readdata),   //                    .readdata
		.out_port   (position28_export)                            // external_connection.export
	);

	nios_system_keycode position_29 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_29_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_29_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_29_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_29_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_29_s1_readdata),   //                    .readdata
		.out_port   (position29_export)                            // external_connection.export
	);

	nios_system_keycode position_3 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_position_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_3_s1_readdata),   //                    .readdata
		.out_port   (position3_export)                            // external_connection.export
	);

	nios_system_keycode position_30 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_30_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_30_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_30_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_30_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_30_s1_readdata),   //                    .readdata
		.out_port   (position30_export)                            // external_connection.export
	);

	nios_system_keycode position_31 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_31_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_31_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_31_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_31_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_31_s1_readdata),   //                    .readdata
		.out_port   (position31_export)                            // external_connection.export
	);

	nios_system_keycode position_32 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_32_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_32_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_32_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_32_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_32_s1_readdata),   //                    .readdata
		.out_port   (position32_export)                            // external_connection.export
	);

	nios_system_keycode position_33 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_33_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_33_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_33_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_33_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_33_s1_readdata),   //                    .readdata
		.out_port   (position33_export)                            // external_connection.export
	);

	nios_system_keycode position_34 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_34_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_34_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_34_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_34_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_34_s1_readdata),   //                    .readdata
		.out_port   (position34_export)                            // external_connection.export
	);

	nios_system_keycode position_35 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_35_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_35_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_35_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_35_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_35_s1_readdata),   //                    .readdata
		.out_port   (position35_export)                            // external_connection.export
	);

	nios_system_keycode position_36 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_position_36_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_36_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_36_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_36_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_36_s1_readdata),   //                    .readdata
		.out_port   (position36_export)                            // external_connection.export
	);

	nios_system_keycode position_4 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_position_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_4_s1_readdata),   //                    .readdata
		.out_port   (position4_export)                            // external_connection.export
	);

	nios_system_keycode position_5 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_position_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_5_s1_readdata),   //                    .readdata
		.out_port   (position5_export)                            // external_connection.export
	);

	nios_system_keycode position_6 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_position_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_6_s1_readdata),   //                    .readdata
		.out_port   (position6_export)                            // external_connection.export
	);

	nios_system_keycode position_7 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_position_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_7_s1_readdata),   //                    .readdata
		.out_port   (position7_export)                            // external_connection.export
	);

	nios_system_keycode position_8 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_position_8_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_8_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_8_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_8_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_8_s1_readdata),   //                    .readdata
		.out_port   (position8_export)                            // external_connection.export
	);

	nios_system_keycode position_9 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_position_9_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_position_9_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_position_9_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_position_9_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_position_9_s1_readdata),   //                    .readdata
		.out_port   (position9_export)                            // external_connection.export
	);

	nios_system_sdram sdram (
		.clk            (sdram_pll_c0_clk),                         //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	nios_system_sdram_pll sdram_pll (
		.clk                (clk_clk),                                         //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),              // inclk_interface_reset.reset
		.read               (mm_interconnect_0_sdram_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_sdram_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_sdram_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_sdram_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_sdram_pll_pll_slave_writedata), //                      .writedata
		.c0                 (sdram_pll_c0_clk),                                //                    c0.clk
		.c1                 (sdram_clk_clk),                                   //                    c1.clk
		.scandone           (),                                                //           (terminated)
		.scandataout        (),                                                //           (terminated)
		.areset             (1'b0),                                            //           (terminated)
		.locked             (),                                                //           (terminated)
		.phasedone          (),                                                //           (terminated)
		.phasecounterselect (4'b0000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                            //           (terminated)
		.phasestep          (1'b0),                                            //           (terminated)
		.scanclk            (1'b0),                                            //           (terminated)
		.scanclkena         (1'b0),                                            //           (terminated)
		.scandata           (1'b0),                                            //           (terminated)
		.configupdate       (1'b0)                                             //           (terminated)
	);

	nios_system_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.sdram_pll_c0_clk                               (sdram_pll_c0_clk),                                            //                             sdram_pll_c0.clk
		.jtag_uart_0_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                              //  jtag_uart_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.sdram_reset_reset_bridge_in_reset_reset        (rst_controller_002_reset_out_reset),                          //        sdram_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.is_new_game_start_s1_address                   (mm_interconnect_0_is_new_game_start_s1_address),              //                     is_new_game_start_s1.address
		.is_new_game_start_s1_readdata                  (mm_interconnect_0_is_new_game_start_s1_readdata),             //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.keycode_s1_address                             (mm_interconnect_0_keycode_s1_address),                        //                               keycode_s1.address
		.keycode_s1_write                               (mm_interconnect_0_keycode_s1_write),                          //                                         .write
		.keycode_s1_readdata                            (mm_interconnect_0_keycode_s1_readdata),                       //                                         .readdata
		.keycode_s1_writedata                           (mm_interconnect_0_keycode_s1_writedata),                      //                                         .writedata
		.keycode_s1_chipselect                          (mm_interconnect_0_keycode_s1_chipselect),                     //                                         .chipselect
		.keycode_0_s1_address                           (mm_interconnect_0_keycode_0_s1_address),                      //                             keycode_0_s1.address
		.keycode_0_s1_write                             (mm_interconnect_0_keycode_0_s1_write),                        //                                         .write
		.keycode_0_s1_readdata                          (mm_interconnect_0_keycode_0_s1_readdata),                     //                                         .readdata
		.keycode_0_s1_writedata                         (mm_interconnect_0_keycode_0_s1_writedata),                    //                                         .writedata
		.keycode_0_s1_chipselect                        (mm_interconnect_0_keycode_0_s1_chipselect),                   //                                         .chipselect
		.keycode_1_s1_address                           (mm_interconnect_0_keycode_1_s1_address),                      //                             keycode_1_s1.address
		.keycode_1_s1_write                             (mm_interconnect_0_keycode_1_s1_write),                        //                                         .write
		.keycode_1_s1_readdata                          (mm_interconnect_0_keycode_1_s1_readdata),                     //                                         .readdata
		.keycode_1_s1_writedata                         (mm_interconnect_0_keycode_1_s1_writedata),                    //                                         .writedata
		.keycode_1_s1_chipselect                        (mm_interconnect_0_keycode_1_s1_chipselect),                   //                                         .chipselect
		.keycode_2_s1_address                           (mm_interconnect_0_keycode_2_s1_address),                      //                             keycode_2_s1.address
		.keycode_2_s1_write                             (mm_interconnect_0_keycode_2_s1_write),                        //                                         .write
		.keycode_2_s1_readdata                          (mm_interconnect_0_keycode_2_s1_readdata),                     //                                         .readdata
		.keycode_2_s1_writedata                         (mm_interconnect_0_keycode_2_s1_writedata),                    //                                         .writedata
		.keycode_2_s1_chipselect                        (mm_interconnect_0_keycode_2_s1_chipselect),                   //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),               //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                         .clken
		.otg_hpi_address_s1_address                     (mm_interconnect_0_otg_hpi_address_s1_address),                //                       otg_hpi_address_s1.address
		.otg_hpi_address_s1_write                       (mm_interconnect_0_otg_hpi_address_s1_write),                  //                                         .write
		.otg_hpi_address_s1_readdata                    (mm_interconnect_0_otg_hpi_address_s1_readdata),               //                                         .readdata
		.otg_hpi_address_s1_writedata                   (mm_interconnect_0_otg_hpi_address_s1_writedata),              //                                         .writedata
		.otg_hpi_address_s1_chipselect                  (mm_interconnect_0_otg_hpi_address_s1_chipselect),             //                                         .chipselect
		.otg_hpi_cs_s1_address                          (mm_interconnect_0_otg_hpi_cs_s1_address),                     //                            otg_hpi_cs_s1.address
		.otg_hpi_cs_s1_write                            (mm_interconnect_0_otg_hpi_cs_s1_write),                       //                                         .write
		.otg_hpi_cs_s1_readdata                         (mm_interconnect_0_otg_hpi_cs_s1_readdata),                    //                                         .readdata
		.otg_hpi_cs_s1_writedata                        (mm_interconnect_0_otg_hpi_cs_s1_writedata),                   //                                         .writedata
		.otg_hpi_cs_s1_chipselect                       (mm_interconnect_0_otg_hpi_cs_s1_chipselect),                  //                                         .chipselect
		.otg_hpi_data_s1_address                        (mm_interconnect_0_otg_hpi_data_s1_address),                   //                          otg_hpi_data_s1.address
		.otg_hpi_data_s1_write                          (mm_interconnect_0_otg_hpi_data_s1_write),                     //                                         .write
		.otg_hpi_data_s1_readdata                       (mm_interconnect_0_otg_hpi_data_s1_readdata),                  //                                         .readdata
		.otg_hpi_data_s1_writedata                      (mm_interconnect_0_otg_hpi_data_s1_writedata),                 //                                         .writedata
		.otg_hpi_data_s1_chipselect                     (mm_interconnect_0_otg_hpi_data_s1_chipselect),                //                                         .chipselect
		.otg_hpi_r_s1_address                           (mm_interconnect_0_otg_hpi_r_s1_address),                      //                             otg_hpi_r_s1.address
		.otg_hpi_r_s1_write                             (mm_interconnect_0_otg_hpi_r_s1_write),                        //                                         .write
		.otg_hpi_r_s1_readdata                          (mm_interconnect_0_otg_hpi_r_s1_readdata),                     //                                         .readdata
		.otg_hpi_r_s1_writedata                         (mm_interconnect_0_otg_hpi_r_s1_writedata),                    //                                         .writedata
		.otg_hpi_r_s1_chipselect                        (mm_interconnect_0_otg_hpi_r_s1_chipselect),                   //                                         .chipselect
		.otg_hpi_reset_s1_address                       (mm_interconnect_0_otg_hpi_reset_s1_address),                  //                         otg_hpi_reset_s1.address
		.otg_hpi_reset_s1_write                         (mm_interconnect_0_otg_hpi_reset_s1_write),                    //                                         .write
		.otg_hpi_reset_s1_readdata                      (mm_interconnect_0_otg_hpi_reset_s1_readdata),                 //                                         .readdata
		.otg_hpi_reset_s1_writedata                     (mm_interconnect_0_otg_hpi_reset_s1_writedata),                //                                         .writedata
		.otg_hpi_reset_s1_chipselect                    (mm_interconnect_0_otg_hpi_reset_s1_chipselect),               //                                         .chipselect
		.otg_hpi_w_s1_address                           (mm_interconnect_0_otg_hpi_w_s1_address),                      //                             otg_hpi_w_s1.address
		.otg_hpi_w_s1_write                             (mm_interconnect_0_otg_hpi_w_s1_write),                        //                                         .write
		.otg_hpi_w_s1_readdata                          (mm_interconnect_0_otg_hpi_w_s1_readdata),                     //                                         .readdata
		.otg_hpi_w_s1_writedata                         (mm_interconnect_0_otg_hpi_w_s1_writedata),                    //                                         .writedata
		.otg_hpi_w_s1_chipselect                        (mm_interconnect_0_otg_hpi_w_s1_chipselect),                   //                                         .chipselect
		.position_0_s1_address                          (mm_interconnect_0_position_0_s1_address),                     //                            position_0_s1.address
		.position_0_s1_write                            (mm_interconnect_0_position_0_s1_write),                       //                                         .write
		.position_0_s1_readdata                         (mm_interconnect_0_position_0_s1_readdata),                    //                                         .readdata
		.position_0_s1_writedata                        (mm_interconnect_0_position_0_s1_writedata),                   //                                         .writedata
		.position_0_s1_chipselect                       (mm_interconnect_0_position_0_s1_chipselect),                  //                                         .chipselect
		.position_1_s1_address                          (mm_interconnect_0_position_1_s1_address),                     //                            position_1_s1.address
		.position_1_s1_write                            (mm_interconnect_0_position_1_s1_write),                       //                                         .write
		.position_1_s1_readdata                         (mm_interconnect_0_position_1_s1_readdata),                    //                                         .readdata
		.position_1_s1_writedata                        (mm_interconnect_0_position_1_s1_writedata),                   //                                         .writedata
		.position_1_s1_chipselect                       (mm_interconnect_0_position_1_s1_chipselect),                  //                                         .chipselect
		.position_10_s1_address                         (mm_interconnect_0_position_10_s1_address),                    //                           position_10_s1.address
		.position_10_s1_write                           (mm_interconnect_0_position_10_s1_write),                      //                                         .write
		.position_10_s1_readdata                        (mm_interconnect_0_position_10_s1_readdata),                   //                                         .readdata
		.position_10_s1_writedata                       (mm_interconnect_0_position_10_s1_writedata),                  //                                         .writedata
		.position_10_s1_chipselect                      (mm_interconnect_0_position_10_s1_chipselect),                 //                                         .chipselect
		.position_11_s1_address                         (mm_interconnect_0_position_11_s1_address),                    //                           position_11_s1.address
		.position_11_s1_write                           (mm_interconnect_0_position_11_s1_write),                      //                                         .write
		.position_11_s1_readdata                        (mm_interconnect_0_position_11_s1_readdata),                   //                                         .readdata
		.position_11_s1_writedata                       (mm_interconnect_0_position_11_s1_writedata),                  //                                         .writedata
		.position_11_s1_chipselect                      (mm_interconnect_0_position_11_s1_chipselect),                 //                                         .chipselect
		.position_12_s1_address                         (mm_interconnect_0_position_12_s1_address),                    //                           position_12_s1.address
		.position_12_s1_write                           (mm_interconnect_0_position_12_s1_write),                      //                                         .write
		.position_12_s1_readdata                        (mm_interconnect_0_position_12_s1_readdata),                   //                                         .readdata
		.position_12_s1_writedata                       (mm_interconnect_0_position_12_s1_writedata),                  //                                         .writedata
		.position_12_s1_chipselect                      (mm_interconnect_0_position_12_s1_chipselect),                 //                                         .chipselect
		.position_13_s1_address                         (mm_interconnect_0_position_13_s1_address),                    //                           position_13_s1.address
		.position_13_s1_write                           (mm_interconnect_0_position_13_s1_write),                      //                                         .write
		.position_13_s1_readdata                        (mm_interconnect_0_position_13_s1_readdata),                   //                                         .readdata
		.position_13_s1_writedata                       (mm_interconnect_0_position_13_s1_writedata),                  //                                         .writedata
		.position_13_s1_chipselect                      (mm_interconnect_0_position_13_s1_chipselect),                 //                                         .chipselect
		.position_14_s1_address                         (mm_interconnect_0_position_14_s1_address),                    //                           position_14_s1.address
		.position_14_s1_write                           (mm_interconnect_0_position_14_s1_write),                      //                                         .write
		.position_14_s1_readdata                        (mm_interconnect_0_position_14_s1_readdata),                   //                                         .readdata
		.position_14_s1_writedata                       (mm_interconnect_0_position_14_s1_writedata),                  //                                         .writedata
		.position_14_s1_chipselect                      (mm_interconnect_0_position_14_s1_chipselect),                 //                                         .chipselect
		.position_15_s1_address                         (mm_interconnect_0_position_15_s1_address),                    //                           position_15_s1.address
		.position_15_s1_write                           (mm_interconnect_0_position_15_s1_write),                      //                                         .write
		.position_15_s1_readdata                        (mm_interconnect_0_position_15_s1_readdata),                   //                                         .readdata
		.position_15_s1_writedata                       (mm_interconnect_0_position_15_s1_writedata),                  //                                         .writedata
		.position_15_s1_chipselect                      (mm_interconnect_0_position_15_s1_chipselect),                 //                                         .chipselect
		.position_16_s1_address                         (mm_interconnect_0_position_16_s1_address),                    //                           position_16_s1.address
		.position_16_s1_write                           (mm_interconnect_0_position_16_s1_write),                      //                                         .write
		.position_16_s1_readdata                        (mm_interconnect_0_position_16_s1_readdata),                   //                                         .readdata
		.position_16_s1_writedata                       (mm_interconnect_0_position_16_s1_writedata),                  //                                         .writedata
		.position_16_s1_chipselect                      (mm_interconnect_0_position_16_s1_chipselect),                 //                                         .chipselect
		.position_17_s1_address                         (mm_interconnect_0_position_17_s1_address),                    //                           position_17_s1.address
		.position_17_s1_write                           (mm_interconnect_0_position_17_s1_write),                      //                                         .write
		.position_17_s1_readdata                        (mm_interconnect_0_position_17_s1_readdata),                   //                                         .readdata
		.position_17_s1_writedata                       (mm_interconnect_0_position_17_s1_writedata),                  //                                         .writedata
		.position_17_s1_chipselect                      (mm_interconnect_0_position_17_s1_chipselect),                 //                                         .chipselect
		.position_18_s1_address                         (mm_interconnect_0_position_18_s1_address),                    //                           position_18_s1.address
		.position_18_s1_write                           (mm_interconnect_0_position_18_s1_write),                      //                                         .write
		.position_18_s1_readdata                        (mm_interconnect_0_position_18_s1_readdata),                   //                                         .readdata
		.position_18_s1_writedata                       (mm_interconnect_0_position_18_s1_writedata),                  //                                         .writedata
		.position_18_s1_chipselect                      (mm_interconnect_0_position_18_s1_chipselect),                 //                                         .chipselect
		.position_19_s1_address                         (mm_interconnect_0_position_19_s1_address),                    //                           position_19_s1.address
		.position_19_s1_write                           (mm_interconnect_0_position_19_s1_write),                      //                                         .write
		.position_19_s1_readdata                        (mm_interconnect_0_position_19_s1_readdata),                   //                                         .readdata
		.position_19_s1_writedata                       (mm_interconnect_0_position_19_s1_writedata),                  //                                         .writedata
		.position_19_s1_chipselect                      (mm_interconnect_0_position_19_s1_chipselect),                 //                                         .chipselect
		.position_2_s1_address                          (mm_interconnect_0_position_2_s1_address),                     //                            position_2_s1.address
		.position_2_s1_write                            (mm_interconnect_0_position_2_s1_write),                       //                                         .write
		.position_2_s1_readdata                         (mm_interconnect_0_position_2_s1_readdata),                    //                                         .readdata
		.position_2_s1_writedata                        (mm_interconnect_0_position_2_s1_writedata),                   //                                         .writedata
		.position_2_s1_chipselect                       (mm_interconnect_0_position_2_s1_chipselect),                  //                                         .chipselect
		.position_20_s1_address                         (mm_interconnect_0_position_20_s1_address),                    //                           position_20_s1.address
		.position_20_s1_write                           (mm_interconnect_0_position_20_s1_write),                      //                                         .write
		.position_20_s1_readdata                        (mm_interconnect_0_position_20_s1_readdata),                   //                                         .readdata
		.position_20_s1_writedata                       (mm_interconnect_0_position_20_s1_writedata),                  //                                         .writedata
		.position_20_s1_chipselect                      (mm_interconnect_0_position_20_s1_chipselect),                 //                                         .chipselect
		.position_21_s1_address                         (mm_interconnect_0_position_21_s1_address),                    //                           position_21_s1.address
		.position_21_s1_write                           (mm_interconnect_0_position_21_s1_write),                      //                                         .write
		.position_21_s1_readdata                        (mm_interconnect_0_position_21_s1_readdata),                   //                                         .readdata
		.position_21_s1_writedata                       (mm_interconnect_0_position_21_s1_writedata),                  //                                         .writedata
		.position_21_s1_chipselect                      (mm_interconnect_0_position_21_s1_chipselect),                 //                                         .chipselect
		.position_22_s1_address                         (mm_interconnect_0_position_22_s1_address),                    //                           position_22_s1.address
		.position_22_s1_write                           (mm_interconnect_0_position_22_s1_write),                      //                                         .write
		.position_22_s1_readdata                        (mm_interconnect_0_position_22_s1_readdata),                   //                                         .readdata
		.position_22_s1_writedata                       (mm_interconnect_0_position_22_s1_writedata),                  //                                         .writedata
		.position_22_s1_chipselect                      (mm_interconnect_0_position_22_s1_chipselect),                 //                                         .chipselect
		.position_23_s1_address                         (mm_interconnect_0_position_23_s1_address),                    //                           position_23_s1.address
		.position_23_s1_write                           (mm_interconnect_0_position_23_s1_write),                      //                                         .write
		.position_23_s1_readdata                        (mm_interconnect_0_position_23_s1_readdata),                   //                                         .readdata
		.position_23_s1_writedata                       (mm_interconnect_0_position_23_s1_writedata),                  //                                         .writedata
		.position_23_s1_chipselect                      (mm_interconnect_0_position_23_s1_chipselect),                 //                                         .chipselect
		.position_24_s1_address                         (mm_interconnect_0_position_24_s1_address),                    //                           position_24_s1.address
		.position_24_s1_write                           (mm_interconnect_0_position_24_s1_write),                      //                                         .write
		.position_24_s1_readdata                        (mm_interconnect_0_position_24_s1_readdata),                   //                                         .readdata
		.position_24_s1_writedata                       (mm_interconnect_0_position_24_s1_writedata),                  //                                         .writedata
		.position_24_s1_chipselect                      (mm_interconnect_0_position_24_s1_chipselect),                 //                                         .chipselect
		.position_25_s1_address                         (mm_interconnect_0_position_25_s1_address),                    //                           position_25_s1.address
		.position_25_s1_write                           (mm_interconnect_0_position_25_s1_write),                      //                                         .write
		.position_25_s1_readdata                        (mm_interconnect_0_position_25_s1_readdata),                   //                                         .readdata
		.position_25_s1_writedata                       (mm_interconnect_0_position_25_s1_writedata),                  //                                         .writedata
		.position_25_s1_chipselect                      (mm_interconnect_0_position_25_s1_chipselect),                 //                                         .chipselect
		.position_26_s1_address                         (mm_interconnect_0_position_26_s1_address),                    //                           position_26_s1.address
		.position_26_s1_write                           (mm_interconnect_0_position_26_s1_write),                      //                                         .write
		.position_26_s1_readdata                        (mm_interconnect_0_position_26_s1_readdata),                   //                                         .readdata
		.position_26_s1_writedata                       (mm_interconnect_0_position_26_s1_writedata),                  //                                         .writedata
		.position_26_s1_chipselect                      (mm_interconnect_0_position_26_s1_chipselect),                 //                                         .chipselect
		.position_27_s1_address                         (mm_interconnect_0_position_27_s1_address),                    //                           position_27_s1.address
		.position_27_s1_write                           (mm_interconnect_0_position_27_s1_write),                      //                                         .write
		.position_27_s1_readdata                        (mm_interconnect_0_position_27_s1_readdata),                   //                                         .readdata
		.position_27_s1_writedata                       (mm_interconnect_0_position_27_s1_writedata),                  //                                         .writedata
		.position_27_s1_chipselect                      (mm_interconnect_0_position_27_s1_chipselect),                 //                                         .chipselect
		.position_28_s1_address                         (mm_interconnect_0_position_28_s1_address),                    //                           position_28_s1.address
		.position_28_s1_write                           (mm_interconnect_0_position_28_s1_write),                      //                                         .write
		.position_28_s1_readdata                        (mm_interconnect_0_position_28_s1_readdata),                   //                                         .readdata
		.position_28_s1_writedata                       (mm_interconnect_0_position_28_s1_writedata),                  //                                         .writedata
		.position_28_s1_chipselect                      (mm_interconnect_0_position_28_s1_chipselect),                 //                                         .chipselect
		.position_29_s1_address                         (mm_interconnect_0_position_29_s1_address),                    //                           position_29_s1.address
		.position_29_s1_write                           (mm_interconnect_0_position_29_s1_write),                      //                                         .write
		.position_29_s1_readdata                        (mm_interconnect_0_position_29_s1_readdata),                   //                                         .readdata
		.position_29_s1_writedata                       (mm_interconnect_0_position_29_s1_writedata),                  //                                         .writedata
		.position_29_s1_chipselect                      (mm_interconnect_0_position_29_s1_chipselect),                 //                                         .chipselect
		.position_3_s1_address                          (mm_interconnect_0_position_3_s1_address),                     //                            position_3_s1.address
		.position_3_s1_write                            (mm_interconnect_0_position_3_s1_write),                       //                                         .write
		.position_3_s1_readdata                         (mm_interconnect_0_position_3_s1_readdata),                    //                                         .readdata
		.position_3_s1_writedata                        (mm_interconnect_0_position_3_s1_writedata),                   //                                         .writedata
		.position_3_s1_chipselect                       (mm_interconnect_0_position_3_s1_chipselect),                  //                                         .chipselect
		.position_30_s1_address                         (mm_interconnect_0_position_30_s1_address),                    //                           position_30_s1.address
		.position_30_s1_write                           (mm_interconnect_0_position_30_s1_write),                      //                                         .write
		.position_30_s1_readdata                        (mm_interconnect_0_position_30_s1_readdata),                   //                                         .readdata
		.position_30_s1_writedata                       (mm_interconnect_0_position_30_s1_writedata),                  //                                         .writedata
		.position_30_s1_chipselect                      (mm_interconnect_0_position_30_s1_chipselect),                 //                                         .chipselect
		.position_31_s1_address                         (mm_interconnect_0_position_31_s1_address),                    //                           position_31_s1.address
		.position_31_s1_write                           (mm_interconnect_0_position_31_s1_write),                      //                                         .write
		.position_31_s1_readdata                        (mm_interconnect_0_position_31_s1_readdata),                   //                                         .readdata
		.position_31_s1_writedata                       (mm_interconnect_0_position_31_s1_writedata),                  //                                         .writedata
		.position_31_s1_chipselect                      (mm_interconnect_0_position_31_s1_chipselect),                 //                                         .chipselect
		.position_32_s1_address                         (mm_interconnect_0_position_32_s1_address),                    //                           position_32_s1.address
		.position_32_s1_write                           (mm_interconnect_0_position_32_s1_write),                      //                                         .write
		.position_32_s1_readdata                        (mm_interconnect_0_position_32_s1_readdata),                   //                                         .readdata
		.position_32_s1_writedata                       (mm_interconnect_0_position_32_s1_writedata),                  //                                         .writedata
		.position_32_s1_chipselect                      (mm_interconnect_0_position_32_s1_chipselect),                 //                                         .chipselect
		.position_33_s1_address                         (mm_interconnect_0_position_33_s1_address),                    //                           position_33_s1.address
		.position_33_s1_write                           (mm_interconnect_0_position_33_s1_write),                      //                                         .write
		.position_33_s1_readdata                        (mm_interconnect_0_position_33_s1_readdata),                   //                                         .readdata
		.position_33_s1_writedata                       (mm_interconnect_0_position_33_s1_writedata),                  //                                         .writedata
		.position_33_s1_chipselect                      (mm_interconnect_0_position_33_s1_chipselect),                 //                                         .chipselect
		.position_34_s1_address                         (mm_interconnect_0_position_34_s1_address),                    //                           position_34_s1.address
		.position_34_s1_write                           (mm_interconnect_0_position_34_s1_write),                      //                                         .write
		.position_34_s1_readdata                        (mm_interconnect_0_position_34_s1_readdata),                   //                                         .readdata
		.position_34_s1_writedata                       (mm_interconnect_0_position_34_s1_writedata),                  //                                         .writedata
		.position_34_s1_chipselect                      (mm_interconnect_0_position_34_s1_chipselect),                 //                                         .chipselect
		.position_35_s1_address                         (mm_interconnect_0_position_35_s1_address),                    //                           position_35_s1.address
		.position_35_s1_write                           (mm_interconnect_0_position_35_s1_write),                      //                                         .write
		.position_35_s1_readdata                        (mm_interconnect_0_position_35_s1_readdata),                   //                                         .readdata
		.position_35_s1_writedata                       (mm_interconnect_0_position_35_s1_writedata),                  //                                         .writedata
		.position_35_s1_chipselect                      (mm_interconnect_0_position_35_s1_chipselect),                 //                                         .chipselect
		.position_36_s1_address                         (mm_interconnect_0_position_36_s1_address),                    //                           position_36_s1.address
		.position_36_s1_write                           (mm_interconnect_0_position_36_s1_write),                      //                                         .write
		.position_36_s1_readdata                        (mm_interconnect_0_position_36_s1_readdata),                   //                                         .readdata
		.position_36_s1_writedata                       (mm_interconnect_0_position_36_s1_writedata),                  //                                         .writedata
		.position_36_s1_chipselect                      (mm_interconnect_0_position_36_s1_chipselect),                 //                                         .chipselect
		.position_4_s1_address                          (mm_interconnect_0_position_4_s1_address),                     //                            position_4_s1.address
		.position_4_s1_write                            (mm_interconnect_0_position_4_s1_write),                       //                                         .write
		.position_4_s1_readdata                         (mm_interconnect_0_position_4_s1_readdata),                    //                                         .readdata
		.position_4_s1_writedata                        (mm_interconnect_0_position_4_s1_writedata),                   //                                         .writedata
		.position_4_s1_chipselect                       (mm_interconnect_0_position_4_s1_chipselect),                  //                                         .chipselect
		.position_5_s1_address                          (mm_interconnect_0_position_5_s1_address),                     //                            position_5_s1.address
		.position_5_s1_write                            (mm_interconnect_0_position_5_s1_write),                       //                                         .write
		.position_5_s1_readdata                         (mm_interconnect_0_position_5_s1_readdata),                    //                                         .readdata
		.position_5_s1_writedata                        (mm_interconnect_0_position_5_s1_writedata),                   //                                         .writedata
		.position_5_s1_chipselect                       (mm_interconnect_0_position_5_s1_chipselect),                  //                                         .chipselect
		.position_6_s1_address                          (mm_interconnect_0_position_6_s1_address),                     //                            position_6_s1.address
		.position_6_s1_write                            (mm_interconnect_0_position_6_s1_write),                       //                                         .write
		.position_6_s1_readdata                         (mm_interconnect_0_position_6_s1_readdata),                    //                                         .readdata
		.position_6_s1_writedata                        (mm_interconnect_0_position_6_s1_writedata),                   //                                         .writedata
		.position_6_s1_chipselect                       (mm_interconnect_0_position_6_s1_chipselect),                  //                                         .chipselect
		.position_7_s1_address                          (mm_interconnect_0_position_7_s1_address),                     //                            position_7_s1.address
		.position_7_s1_write                            (mm_interconnect_0_position_7_s1_write),                       //                                         .write
		.position_7_s1_readdata                         (mm_interconnect_0_position_7_s1_readdata),                    //                                         .readdata
		.position_7_s1_writedata                        (mm_interconnect_0_position_7_s1_writedata),                   //                                         .writedata
		.position_7_s1_chipselect                       (mm_interconnect_0_position_7_s1_chipselect),                  //                                         .chipselect
		.position_8_s1_address                          (mm_interconnect_0_position_8_s1_address),                     //                            position_8_s1.address
		.position_8_s1_write                            (mm_interconnect_0_position_8_s1_write),                       //                                         .write
		.position_8_s1_readdata                         (mm_interconnect_0_position_8_s1_readdata),                    //                                         .readdata
		.position_8_s1_writedata                        (mm_interconnect_0_position_8_s1_writedata),                   //                                         .writedata
		.position_8_s1_chipselect                       (mm_interconnect_0_position_8_s1_chipselect),                  //                                         .chipselect
		.position_9_s1_address                          (mm_interconnect_0_position_9_s1_address),                     //                            position_9_s1.address
		.position_9_s1_write                            (mm_interconnect_0_position_9_s1_write),                       //                                         .write
		.position_9_s1_readdata                         (mm_interconnect_0_position_9_s1_readdata),                    //                                         .readdata
		.position_9_s1_writedata                        (mm_interconnect_0_position_9_s1_writedata),                   //                                         .writedata
		.position_9_s1_chipselect                       (mm_interconnect_0_position_9_s1_chipselect),                  //                                         .chipselect
		.sdram_s1_address                               (mm_interconnect_0_sdram_s1_address),                          //                                 sdram_s1.address
		.sdram_s1_write                                 (mm_interconnect_0_sdram_s1_write),                            //                                         .write
		.sdram_s1_read                                  (mm_interconnect_0_sdram_s1_read),                             //                                         .read
		.sdram_s1_readdata                              (mm_interconnect_0_sdram_s1_readdata),                         //                                         .readdata
		.sdram_s1_writedata                             (mm_interconnect_0_sdram_s1_writedata),                        //                                         .writedata
		.sdram_s1_byteenable                            (mm_interconnect_0_sdram_s1_byteenable),                       //                                         .byteenable
		.sdram_s1_readdatavalid                         (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                         .readdatavalid
		.sdram_s1_waitrequest                           (mm_interconnect_0_sdram_s1_waitrequest),                      //                                         .waitrequest
		.sdram_s1_chipselect                            (mm_interconnect_0_sdram_s1_chipselect),                       //                                         .chipselect
		.sdram_pll_pll_slave_address                    (mm_interconnect_0_sdram_pll_pll_slave_address),               //                      sdram_pll_pll_slave.address
		.sdram_pll_pll_slave_write                      (mm_interconnect_0_sdram_pll_pll_slave_write),                 //                                         .write
		.sdram_pll_pll_slave_read                       (mm_interconnect_0_sdram_pll_pll_slave_read),                  //                                         .read
		.sdram_pll_pll_slave_readdata                   (mm_interconnect_0_sdram_pll_pll_slave_readdata),              //                                         .readdata
		.sdram_pll_pll_slave_writedata                  (mm_interconnect_0_sdram_pll_pll_slave_writedata),             //                                         .writedata
		.sysid_qsys_0_control_slave_address             (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata            (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)        //                                         .readdata
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (sdram_pll_c0_clk),                       //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
